module hello

pub fn hello() {
	println("Hello World!")
}
